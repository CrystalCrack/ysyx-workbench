`define SINGLE_CYCLE
