module LSU(

);

endmodule
