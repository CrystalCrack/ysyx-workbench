// `define CONFIG_DSTAGE_BUF
`define CONFIG_XSTAGE_BUF
`define CONFIG_MSTAGE_BUF
`define CONFIG_WSTAGE_BUF






